//Ethan Sarif-Kattan & LH Lee

package uart_tx_pkg;
    `include "uart_tx_transaction.sv"
    `include "uart_tx_generator.sv"
    `include "uart_tx_driver.sv"
    `include "uart_tx_monitor.sv"
    `include "uart_tx_scoreboard.sv"
    `include "uart_tx_environment.sv"
    `include "uart_tx_test.sv" 
 
endpackage : uart_tx_pkg

// `include "interface.sv"

