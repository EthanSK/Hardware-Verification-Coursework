package ahb_uart_pkg;
    `include "ahb_uart_transaction.sv"
    `include "ahb_uart_generator.sv"
    `include "ahb_uart_tx_driver.sv"
    `include "ahb_uart_tx_monitor.sv"
    `include "ahb_uart_tx_scoreboard.sv"
    `include "ahb_uart_environment.sv"
    `include "ahb_uart_test.sv" 
 
endpackage : ahb_uart_pkg

// `include "interface.sv"

