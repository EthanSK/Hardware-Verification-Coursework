class transaction;

    rand bit [8:0] d_in;
    bit [8:0] d_out;
 
endclass