package uart_rx_pkg;
    `include "uart_rx_transaction.sv"
    `include "uart_rx_generator.sv"
    `include "uart_rx_driver.sv"
    `include "uart_rx_monitor.sv"
    `include "uart_rx_scoreboard.sv"
    `include "uart_rx_environment.sv"
    `include "uart_rx_test.sv" 
 
endpackage : uart_rx_pkg

// `include "interface.sv"

