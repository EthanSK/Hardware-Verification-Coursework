package parity_check_pkg;
    `include "parity_check_transaction.sv"
    `include "parity_check_generator.sv"
    `include "parity_check_runner.sv"
    `include "parity_check_scoreboard.sv"
    `include "parity_check_environment.sv"
    `include "parity_check_test.sv" 

endpackage : parity_check_pkg

