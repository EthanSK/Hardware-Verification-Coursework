import pkg:test;

module testbench;
    reg clk;
    reg baud_tick;

    _if _if(clk, baud_tick);

    

    initial begin
        
    end
endmodule