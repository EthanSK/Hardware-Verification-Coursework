//Ethan Sarif-Kattan & LH Lee

package ahblite_sys_pkg;
    `include "ahblite_sys_transaction.sv"
    `include "ahblite_sys_generator.sv"
    `include "ahblite_sys_driver.sv"
    `include "ahblite_sys_monitor.sv"
    `include "ahblite_sys_scoreboard.sv"
    `include "ahblite_sys_environment.sv"
    `include "ahblite_sys_test.sv" 
 
endpackage : ahblite_sys_pkg

