package pkg;
    `include "driver.sv"
    `include "environment.sv"
    `include "monitor.sv"
    `include "scoreboard.sv"
    `include "test.sv"
    `include "transaction.sv"
endpackage : pkg

    `include "interface.sv"